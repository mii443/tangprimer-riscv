`define OP_SW      32'b00000000000000000010000000100011
`define MASK_OP_SW 32'b00000000000000000111000001111111

`define OP_LW      32'b00000000000000000010000000000011
`define MASK_OP_LW 32'b00000000000000000111000001111111

`define OP_LUI      32'b00000000000000000000000000110111
`define MASK_OP_LUI 32'b00000000000000000000000001111111

`define OP_ADDI      32'b00000000000000000000000000010011
`define MASK_OP_ADDI 32'b00000000000000000111000001111111