`define OP_SW 7'b0100011
`define OP_LW 7'b0000011